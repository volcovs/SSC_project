library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;


entity HardDisk is
    port (clk: in STD_LOGIC;
        enable: in STD_LOGIC;
        write: in STD_LOGIC;
        -- adresa contine numarul paginii fizice si offset-ul la care se gaseste cuvantul de citit
        -- 18 biti => numarul paginii, 12 biti => offset-ul (daca octeti individuali)
        -- scaled down => 5 biti/pagina, 4 biti/offset
        read_address: in STD_LOGIC_VECTOR(8 downto 0);
        write_address: in STD_LOGIC_VECTOR(8 downto 0);
        -- magistrala de date este pe 16 biti, de aceea blocul de scriere/citire e tot de 16 biti
        WriteData: in STD_LOGIC_VECTOR(15 downto 0);
        ReadData: out STD_LOGIC_VECTOR(15 downto 0));
end HardDisk;

architecture Behavioral of HardDisk is

-- o pagina are 4KB de date => 4096 de bytes
-- scaled down => pagina de 128 de biti
type page is array (0 to 2**4-1) of STD_LOGIC_VECTOR(7 downto 0);
-- intreaga memorie are 2^18 de pagini
-- scaled down => 32 de pagini
type mem is array (0 to 31) of page;

signal pageNumRead: STD_LOGIC_VECTOR(4 downto 0);
signal pageOffsetRead: STD_LOGIC_VECTOR(3 downto 0);
signal pageNumWrite: STD_LOGIC_VECTOR(4 downto 0);
signal pageOffsetWrite: STD_LOGIC_VECTOR(3 downto 0);    

signal memory: mem := (
    -- page 0
    ("10111001", "01100110", "11001001", "00111101",
    "11100010", "01011000", "10010110", "00101001",
    "11000101", "10110101", "00010011", "11100101",
    "01011011", "11100100", "00101011", "10001110"),
    
    -- page 1
    ("11100101", "01010110", "10011001", "00110101",
    "11001010", "01101100", "10100101", "00011101",
    "11101001", "10010101", "00110011", "11001101",
    "01011001", "10110100", "00011011", "11101100"),
    
    -- page 2
    ("10101100", "01101010", "11011001", "00111100",
    "11100110", "01001001", "10010111", "00100011",
    "11001101", "10111101", "00011110", "11101001",
    "01010110", "10101001", "00111001", "11000111"),
    
    -- page 3
    ("11011010", "01001110", "11100101", "00110110",
    "10101001", "01111101", "10010100", "00100011",
    "11100111", "10011001", "01001101", "10110101",
    "00011010", "11101001", "01010110", "10101101"),
    
    -- page 4 
    ("00010001", "00001110", "00000011", "00000100",
    "00000101", "00000110", "00000111", "00001000",
    "00001001", "00001010", "00001011", "00001100",
    "00001101", "00001110", "00001111", "00010000"),
    
    -- page 5
    ("01101010", "00111001", "11000101", "01001111",     
    "10101010", "11110001", "00010101", "10011001",
    "01101000", "10111011", "00111110", "01000100",
    "11111100", "11001010", "00110101", "10101011"),
    
    -- page 6
    ("10101010", "11001100", "00110011", "11110000",
    "01010101", "00110011", "11111100", "00001111",
    "11100000", "00111100", "11001100", "00001111",
    "00111100", "10101010", "11001100", "01010101"),
    
    -- page 7
    ("11011001", "00110110", "11101001", "01011101",
    "00100010", "10101100", "01111010", "11001001",
    "01001100", "11110101", "10010100", "00111011",
    "01101011", "10011110", "00001101", "11101000"),
    
    -- page 8
    ("00000000", "00000001", "00000010", "00000011",
    "00000100", "00000101", "00000110", "00000111",
    "00001000", "00001001", "00001010", "00000011", 
    "00001100", "00001101", "00001110", "00001111"),
    
    -- page 9 
    ("11001001", "01100110", "10111001", "00101001",
    "11100101", "00010011", "01011011", "00111101",
    "00100110", "10100011", "01110100", "11011011",
    "11101010", "01111011", "10001110", "00011110"),
    
    -- page 10
    ("11001001", "01100110", "10111001", "00101001",
    "11100101", "00010011", "01011011", "00111101",
    "00100110", "10100011", "01110100", "11011011",
    "11101010", "01111011", "10001110", "00011110"),
    
    -- page 11
    ("10111001", "01100110", "11001001", "00111101",
    "11100010", "01011000", "10010110", "00101001",
    "11000101", "10110101", "00010011", "11100101",
    "01011011", "11100100", "00101011", "10001110"),
    
    -- page 12
    ("10111001", "01100110", "11001001", "00111101",
    "11100010", "01011000", "10010110", "00101001",
    "11000101", "10110101", "00010011", "11100101",
    "01011011", "11100100", "00101011", "10001110"),
    
    -- page 13
    ("11001001", "01100110", "10111001", "00101001",
    "11100101", "00010011", "01011011", "00111101",
    "00100110", "10100011", "01110100", "11011011",
    "11101010", "01111011", "10001110", "00011110"),
    
    -- page 14
    ("10111001", "01100110", "11001001", "00111101",
    "11100010", "01011000", "10010110", "00101001",
    "11000101", "10110101", "00010011", "11100101",
    "01011011", "11100100", "00101011", "10001110"),
    
    -- page 15
    ("11001001", "01100110", "10111001", "00101001",
    "11100101", "00010011", "01011011", "00111101",
    "00100110", "10100011", "01110100", "11011011",
    "11101010", "01111011", "10001110", "00011110"),
    
    -- page 16
    ("10111001", "01100110", "11001001", "00111101",
    "11100010", "01011000", "10010110", "00101001",
    "11000101", "10110101", "00010011", "11100101",
    "01011011", "11100100", "00101011", "10001110"),
    
    -- page 17
    ("11001001", "01100110", "10111001", "00101001",
    "11100101", "00010011", "01011011", "00111101",
    "00100110", "10100011", "01110100", "11011011",
    "11101010", "01111011", "10001110", "00011110"),
    
    others => (others => (others => '0')));

begin

    pageNumRead <= read_address(8 downto 4);
    pageOffsetRead <= read_address(3 downto 0);
    pageNumWrite <= write_address(8 downto 4);
    pageOffsetWrite <= write_address(3 downto 0);
    
    
    -- scriere sincrona in memorie
    WRITE_PROC: process(clk, write, enable, WriteData, pageNumWrite, pageOffsetWrite) 
    begin
        if (clk'event and clk = '1') then
            if (write = '1' and enable = '1') then
                memory(conv_integer(pageNumWrite))(conv_integer(pageOffsetWrite)) <= WriteData(7 downto 0);
                memory(conv_integer(pageNumWrite))(conv_integer(pageOffsetWrite)+1) <= WriteData(15 downto 8);
            end if;
        end if;    
    end process;
    
    
    -- citire asincrona din memorie
    ReadData(7 downto 0) <= memory(conv_integer(pageNumRead))(conv_integer(pageOffsetRead));
    ReadData(15 downto 8) <= memory(conv_integer(pageNumRead))(conv_integer(pageOffsetRead)+1);


end Behavioral;
